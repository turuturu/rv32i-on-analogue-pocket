

module alu (
    input logic [31:0] op1,
    input logic [31:0] op2,
    output logic [31:0] result,
    output logic is_branch
);

endmodule